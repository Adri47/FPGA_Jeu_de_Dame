----------------------------------------------------------------------------------
-- Company: ENSEIRB-MATMECA
-- Engineer: Adrien CLAIN
-- 
-- Create Date: 12.03.2021 08:41:06
-- Module Name: affichage_jeu_de_dame - Behavioral
-- Project Name: Jeu de dame
-- Target Devices: Nexys 4

-----------------------------------------------------------------------------------------------
--------------------------- Bloc qui vient lire la m�moire afin de mettre ---------------------
--------------------------- � jour l'affichage du jeu de dame----------------------------------
-----------------------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity affichage_jeu_de_dame is
  Port ( clk                     : in std_logic; 
         rst                     : in std_logic;
         e_affichage_jeu_de_dame : in std_logic;                          -- activation du bloc par la FSM
         e_plateau               : in std_logic_vector(7 downto 0);       -- case m�moire 0 � 99 envoy� par la mem
         s_fin_affichage         : out std_logic;                         -- sortie � 1 d�s que le bloc a termin� l'affichage
         s_data_write            : out std_logic;                         -- activation �criture dans le bloc VGA
         s_RW_mem                : out std_logic;                         -- lecture/ecriture de la m�moire
         s_activation_memoire    : out std_logic;                         -- activation de la R/W de la m�moire
         s_addr_vga              : out std_logic_vector (16 downto 0);    -- addresse du pixel � afficher envoy� au VGA 
         s_plateau               : out std_logic_vector(7 downto 0);      -- choix de la case m�moire � lire dans la mem
         s_data_in               : out std_logic_vector (11 downto 0)     -- donn�e � envoyer au bloc VGA
         );
end affichage_jeu_de_dame;

architecture Behavioral of affichage_jeu_de_dame is

-- Creation de type tableau de 576 cases d'entier qui repr�sente la memoire d'un bloc de 24x24 pixels
TYPE mem_bloc IS ARRAY(0 TO 575) OF integer;   

SIGNAL case_blanche           : mem_bloc := (4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095);
SIGNAL case_noire             : mem_bloc := (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0);
SIGNAL pion_blanc             : mem_bloc := (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0);
SIGNAL pion_marron            : mem_bloc := (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0);
SIGNAL dame_marron            : mem_bloc := (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 0, 0, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 0, 0, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 0, 0, 2096, 2096, 2096, 0, 0, 2096, 0, 2096, 0, 2096, 2096, 2096, 2096, 0, 2096, 0, 2096, 0, 0, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0);
SIGNAL dame_blanche           : mem_bloc := (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 0, 0, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 0, 0, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 0, 0, 4095, 4095, 4095, 0, 0, 4095, 0, 4095, 0, 4095, 4095, 4095, 4095, 0, 4095, 0, 4095, 0, 0, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0);
SIGNAL selection_case_noire   : mem_bloc := (2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816);
SIGNAL selection_case_blanche : mem_bloc := (2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816);
SIGNAL selection_pion_marron  : mem_bloc := (2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 2816, 2816, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2816, 2816, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2816, 2816, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2816, 2816, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2816, 2816, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2816, 2816, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816);
SIGNAL selection_pion_blanc   : mem_bloc := (2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 2816, 2816, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 2816, 2816, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 2816, 2816, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 2816, 2816, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 2816, 2816, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 2816, 2816, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816);
SIGNAL selection_dame_blanche : mem_bloc := (2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 2816, 2816, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 2816, 2816, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 2816, 2816, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 4095, 4095, 0, 0, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 2816, 2816, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 0, 0, 4095, 0, 4095, 0, 4095, 4095, 4095, 4095, 0, 4095, 0, 4095, 0, 0, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 0, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 2816, 2816, 0, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 0, 2816, 2816, 0, 0, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 0, 0, 2816, 2816, 0, 0, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 4095, 0, 4095, 4095, 4095, 4095, 4095, 0, 0, 2816, 2816, 0, 0, 0, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 4095, 0, 0, 0, 0, 0, 0, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816);
SIGNAL selection_dame_marron  : mem_bloc := (2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 2816, 2816, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2816, 2816, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 2816, 2816, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2096, 2096, 0, 0, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2816, 2816, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 0, 0, 2096, 0, 2096, 0, 2096, 2096, 2096, 2096, 0, 2096, 0, 2096, 0, 0, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2816, 2816, 0, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2816, 2816, 0, 0, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 0, 0, 2816, 2816, 0, 0, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 2096, 0, 2096, 2096, 2096, 2096, 2096, 0, 0, 2816, 2816, 0, 0, 0, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 2816, 2816, 0, 0, 0, 0, 0, 0, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 2096, 0, 0, 0, 0, 0, 0, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816, 2816);

SIGNAL buffer_bloc            : mem_bloc;

--Tableau regroupant la liste des premieres addresses pixels de chaque case
TYPE premier_pixel IS ARRAY (0 to 99) of integer;
SIGNAL addr_premier_pixel : premier_pixel := (39, 63, 87, 111, 135, 159, 183, 207, 231, 255, 7719, 7743, 7767, 7791, 7815, 7839, 7863, 7887, 7911, 7935, 15399, 15423, 15447, 15471, 15495, 15519, 15543, 15567, 15591, 15615, 23079, 23103, 23127, 23151, 23175, 23199, 23223, 23247, 23271, 23295, 30759, 30783, 30807, 30831, 30855, 30879, 30903, 30927, 30951, 30975, 38439, 38463, 38487, 38511, 38535, 38559, 38583, 38607, 38631, 38655, 46119, 46143, 46167, 46191, 46215, 46239, 46263, 46287, 46311, 46335, 53799, 53823, 53847, 53871, 53895, 53919, 53943, 53967, 53991, 54015, 61479, 61503, 61527, 61551, 61575, 61599, 61623, 61647, 61671, 61695, 69159, 69183, 69207, 69231, 69255, 69279, 69303, 69327, 69351, 69375);

-- d�claration des �tats de la FSM
TYPE state IS (etatInit, etat1, etat2, etat3, etat4, etat5, etat6, etat7, etat8, etat9, etat10); 
SIGNAL next_state, current_state : state;

signal addr_case_plateau           : integer range 0 to 99;         -- signal representant l'addresse de la case du plateau (plateau = 10 x 10 = 100 blocs avec addr = 0 � 99)
signal activation_cpt_addr_plateau : std_logic;                     -- autorisation d'incrementer addr_plateau
signal fin_ecriture_bloc           : std_logic;                     -- signal activer lors de la fin de l'�criture d'un bloc par le module
signal rst_addr_plateau            : std_logic;                     -- signal de remise � z�ro du compteur d'adresse du plateau
signal activer_ecriture_vga        : std_logic;                     -- signal d'activation du compteur de pixel pour �crire sur le bloc VGA
signal affectation_cpt_addr_pixel  : std_logic;                     -- signal qui permet la recopie du premier pixel dans le compteur

signal buffer_plateau              : std_logic_vector (7 downto 0); -- signal tampon stockant la valeur contenu dans un case m�moire du plateau (de x"00" � x"0b")
signal buff_addr_premier_pixel     : unsigned(16 downto 0);         -- signal tampon stockant l'adresse du premier pixel d'un bloc
signal envoi_data                  : std_logic;
--signaux compteur 
signal cpt                         : unsigned(16 downto 0) := (others => '0'); -- compteur 
signal indice_affichage            : unsigned(9 downto 0)  := (others => '0'); -- compteur parcourant le bloc memoire associ� (0 � 575)
signal y                           : unsigned(4 downto 0)  := (others => '0'); -- nombre de ligne axe Y (0 � 23)
signal cpt_max                     : unsigned(16 downto 0) := (others => '0'); -- max = 320*240 = 76800

begin

-- Compteur des adresses pixels piloter par la FSM
     process(clk, rst) is  
        begin
            if rst = '1' then
                cpt <= (others => '0'); 
                y <= (others => '0');
                indice_affichage <= (others => '0');
                fin_ecriture_bloc <= '0';
                cpt_max <= (others => '0');
                cpt <= (others => '0');
                
            elsif clk'event and clk = '1' then
                if affectation_cpt_addr_pixel = '1' then        --on passe � cette condition si on passe � un new bloc
                    cpt <= buff_addr_premier_pixel;             -- affectation du du new premier pixel
                    fin_ecriture_bloc <= '0';                   -- condition � mettre pour enclencher le cpt
                    indice_affichage <= (others => '0');
                    y <= (others => '0');
                    cpt_max <= (buff_addr_premier_pixel + 23);
                 else
                    if activer_ecriture_vga = '1' then
                        if (y < 24 and fin_ecriture_bloc = '0' and indice_affichage /= 575) then --si on est pas sur la derni�re ligne / si cn a pas fini d'afficher le bloc et si on a pas lu last case m�moire du bloc
                            if (cpt < cpt_max) then
                                cpt <= cpt + 1;
                                indice_affichage <= indice_affichage + 1;
                             elsif cpt < (buff_addr_premier_pixel + 7422) then --320*23+23+39 (dernier pixel en bas � droite)
                                y <= y + 1;                                    -- saut de ligne
                                cpt_max <= cpt_max + 320;                      -- new cpt_ligne � chauqe saut de ligne Y                         
                                cpt <= cpt + 297;                              -- new cpt � chauqe saut de ligne Y (= 320 - 23)
                                indice_affichage <= indice_affichage + 1;     
                             else
                                y <= y + 1;
                             end if;
                          else
                            fin_ecriture_bloc <= '1';
                            y <= (others => '0');                 
                          end if;
                     end if;
                 end if;          
            end if;
        end process;

    process (clk, rst, envoi_data)
        begin
            if rst ='1' then
                  s_addr_vga <= (others => '0');
                  s_data_write <= '0';
                  s_data_in <= (others => '0');
            elsif clk'event and clk = '1' then
                if envoi_data = '1' then
                    s_addr_vga <= std_logic_vector(cpt);
                    s_data_write <= '1';
                    s_data_in <= std_logic_vector(to_unsigned((buffer_bloc(to_integer(indice_affichage))),12));
                end if;
            end if;
        end process;
    
    --  Compteur adresse du plateau (0 � 99)
    process(clk, rst) is  
    begin
        IF rst = '1' THEN
            addr_case_plateau <= 0;
        ELSIF clk'event AND clk = '1' THEN
            if activation_cpt_addr_plateau = '1' then
                addr_case_plateau <= addr_case_plateau + 1;
            elsif rst_addr_plateau = '1' then
                addr_case_plateau <= 0;
            end if;
       END IF;
    end process;
   
-----  FSM de la partie affichage -------
     process (clk, rst) is 
         begin   
           if rst = '1' then
               current_state <= etatInit;
           elsif clk'event and clk = '1' then
                   current_state <= next_state;  
           end if;
     end process;
     
     process(current_state, e_affichage_jeu_de_dame, fin_ecriture_bloc, e_plateau,addr_case_plateau)
        begin
            case current_state is
                when etatInit => 
                    if (e_affichage_jeu_de_dame = '1') then
                        next_state <= etat1;
                    else 
                        next_state <= etatInit;
                    end if;
                
                when etat1 =>
                    next_state <= etat2;
                    
                when etat2 =>
                    next_state <= etat3;
                    
                when etat3 =>
                    next_state <= etat4;
                    
                when etat4 =>
                    next_state <= etat5;
                    
                when etat5 =>
                    next_state <= etat6;
                    
                when etat6 =>
                    next_state <= etat7;
                    
                when etat7 =>
                    if fin_ecriture_bloc = '1' then
                        if addr_case_plateau < 99 then
                            next_state <= etat8;
                        else
                            next_state <= etat9;
                        end if;
                     else
                        next_state <= etat7;
                     end if;   
                                      
                when etat8 =>
                    next_state <= etat1;
                --non utilis� d�sormais mais on garde au cas o�    
                when etat9 =>
                    next_state <= etat10;
                  --non utilis� d�sormais mais on garde au cas o�   
                when etat10 =>
                    next_state <= etatInit;
                                   
            end case;
     end process;

    process(current_state, addr_case_plateau, e_plateau, buffer_plateau,
            case_blanche, case_noire, 
            pion_marron, dame_marron, 
            pion_blanc, dame_blanche, 
            selection_case_blanche, 
            selection_case_noire, 
            selection_dame_marron, 
            selection_pion_blanc, 
            selection_dame_blanche,
            selection_pion_marron)
            
        begin
            case current_state is
            
                when etatInit =>
                --remise � z�ro du cpt des cases m�moire (0 � 99) et activation de la m�moire
                rst_addr_plateau               <= '1'; 
                activer_ecriture_vga           <= '0';
                affectation_cpt_addr_pixel     <= '0';
                activation_cpt_addr_plateau    <= '0';
                s_RW_mem                       <= '0';
                s_activation_memoire           <= '1';  
                s_fin_affichage                <= '0';
                envoi_data                     <= '0';
                s_plateau                      <= (others =>'0');
                buffer_plateau                 <= (others =>'0');
                buff_addr_premier_pixel        <= (others => '0');
                
                when etat1 =>
                    --on demande la lecture de la case m�moire � l'addresse "addr_case_plateau" et on enl�ve la remise � z�ro du compteur d'adresse du plateau
                    s_plateau                   <= std_logic_vector(to_unsigned(addr_case_plateau,8));                        
                    
                    rst_addr_plateau               <= '0'; 
                    activer_ecriture_vga           <= '0';
                    affectation_cpt_addr_pixel     <= '0';
                    activation_cpt_addr_plateau    <= '0';
                    s_RW_mem                       <= '0';
                    s_activation_memoire           <= '1';  
                    s_fin_affichage                <= '0';
                    envoi_data                     <= '0';
                    buffer_plateau                 <= (others =>'0');         
                    buff_addr_premier_pixel        <= (others => '0');
                    
                when etat2 =>
                    --on vient stocker la donn�es envoy�e par la m�moire
                    buffer_plateau <= e_plateau; 
                    
                    rst_addr_plateau               <= '0'; 
                    activer_ecriture_vga           <= '0';
                    affectation_cpt_addr_pixel     <= '0';
                    activation_cpt_addr_plateau    <= '0';
                    s_RW_mem                       <= '0';
                    s_activation_memoire           <= '1';  
                    s_fin_affichage                <= '0';
                    envoi_data                     <= '0';
                    s_plateau                      <= std_logic_vector(to_unsigned(addr_case_plateau,8));
                    buff_addr_premier_pixel        <= (others => '0');
                    
                when etat3 =>
                    -- on affecte dans un buffer la memoire d'un bloc d�termin� par sa valeur stock�e dans buffer_plateau
                    rst_addr_plateau               <= '0'; 
                    activer_ecriture_vga           <= '0';
                    affectation_cpt_addr_pixel     <= '0';
                    activation_cpt_addr_plateau    <= '0';
                    s_RW_mem                       <= '0';
                    s_activation_memoire           <= '0';  
                    s_fin_affichage                <= '0';
                    envoi_data                     <= '0';
                    s_plateau                      <= (others =>'0');
                   -- buffer_plateau                 <= e_plateau;
                    buff_addr_premier_pixel        <= (others => '0');
                   
                    case buffer_plateau is
                    
                        when x"00" =>
                            buffer_bloc <= case_blanche;
                
                        when x"01" =>
                            buffer_bloc <= case_noire;
                            
                        when x"02" =>
                            buffer_bloc <= pion_marron;
                            
                        when x"03" =>
                            buffer_bloc <= dame_marron;
                            
                        when x"04" =>
                            buffer_bloc <= pion_blanc;
                            
                        when x"05" =>
                            buffer_bloc <= dame_blanche;
                            
                        when x"06" =>
                            buffer_bloc <= selection_case_blanche;
                            
                        when x"07" =>
                            buffer_bloc <= selection_case_noire;
                            
                        when x"08" =>
                            buffer_bloc <= selection_pion_marron;
                            
                        when x"09" =>
                            buffer_bloc <= selection_dame_marron;
                            
                        when x"0a" =>
                            buffer_bloc <= selection_pion_blanc;
                            
                        when x"0b" =>
                            buffer_bloc <= selection_dame_blanche;
                        
                        -- faire l'export matlab si le besoin est.
--                        when x"0c" =>
--                            buffer_bloc <=
--                        when x"0d" =>
--                            buffer_bloc <=
                        when others =>
                            buffer_bloc <= selection_dame_marron;
                   end case;
                   
                when etat4 =>
                    -- on affecte dans un buffer le premier pixel correspondant � un bloc qui est stock� dans le tableau "addr_premier_pixel"
                    buff_addr_premier_pixel        <= to_unsigned(addr_premier_pixel(addr_case_plateau),17);
                    
                    rst_addr_plateau               <= '0'; 
                    activer_ecriture_vga           <= '0';
                    affectation_cpt_addr_pixel     <= '0';
                    activation_cpt_addr_plateau    <= '0';
                    s_RW_mem                       <= '0';
                    s_activation_memoire           <= '0';  
                    s_fin_affichage                <= '0';
                    envoi_data                     <= '0';
                    s_plateau                      <= (others =>'0');
                    buffer_plateau                 <= (others =>'0');
                    buff_addr_premier_pixel        <= (others => '0');
                    
                when etat5 =>
                    -- permet d'activer la recopie du premier pixel dans le compteur
                    
                    rst_addr_plateau               <= '0'; 
                    activer_ecriture_vga           <= '0';
                    affectation_cpt_addr_pixel     <= '1';
                    activation_cpt_addr_plateau    <= '0';
                    s_RW_mem                       <= '0';
                    s_activation_memoire           <= '0';  
                    s_fin_affichage                <= '0';
                    envoi_data                     <= '0';
                    s_plateau                      <= (others =>'0');
                    buffer_plateau                 <= (others =>'0');
                    buff_addr_premier_pixel        <= to_unsigned(addr_premier_pixel(addr_case_plateau),17);
                    
                when etat6 =>
                    -- d�sactivation de la recopie

                    rst_addr_plateau               <= '0'; 
                    activer_ecriture_vga           <= '0';
                    affectation_cpt_addr_pixel     <= '0';
                    activation_cpt_addr_plateau    <= '0';
                    s_RW_mem                       <= '0';
                    s_activation_memoire           <= '0';  
                    s_fin_affichage                <= '0';
                    envoi_data                     <= '0';
                    s_plateau                      <= (others =>'0');
                    buffer_plateau                 <= (others =>'0');
                    buff_addr_premier_pixel        <= to_unsigned(addr_premier_pixel(addr_case_plateau),17);
                    
                when etat7 =>
                    -- activation de l'envoie des donn�es au bloc VGA + incr�mentation du cpt adresse VGA

                    rst_addr_plateau               <= '0'; 
                    activer_ecriture_vga           <= '1';
                    affectation_cpt_addr_pixel     <= '0';
                    activation_cpt_addr_plateau    <= '0';
                    s_RW_mem                       <= '0';
                    s_activation_memoire           <= '0';  
                    s_fin_affichage                <= '0';  
                    envoi_data                     <= '1';                    
                    s_plateau                      <= (others =>'0');
                    buffer_plateau                 <= (others =>'0');
                    buff_addr_premier_pixel        <= to_unsigned(addr_premier_pixel(addr_case_plateau),17);
                                     
                when etat8 =>
                    -- d�sactivation de l'envoie des donn�es au bloc VGA + arr�t du cpt adresse + incr�mentation du ctp d'adresse plateau + r�cup�ration du premier pixel du nouveau bloc
                    
                    rst_addr_plateau               <= '0'; 
                    activer_ecriture_vga           <= '0';
                    affectation_cpt_addr_pixel     <= '0';
                    activation_cpt_addr_plateau    <= '1';
                    s_RW_mem                       <= '0';
                    s_activation_memoire           <= '0';  
                    s_fin_affichage                <= '0';
                    envoi_data                     <= '0';
                    s_plateau                      <= (others =>'0');
                    buffer_plateau                 <= (others =>'0');
                    buff_addr_premier_pixel        <= (others => '0');
                --non utilis� d�sormais mais on garde au cas o�     
                when etat9 =>
                    -- on arr�te l'incr�mentation d�s qu'on arrive � la fin du plateau soit � l'addr 99
                    
                    rst_addr_plateau               <= '0'; 
                    activer_ecriture_vga           <= '0';
                    affectation_cpt_addr_pixel     <= '0';
                    activation_cpt_addr_plateau    <= '0';
                    s_RW_mem                       <= '0';
                    s_activation_memoire           <= '0';  
                    s_fin_affichage                <= '0';
                    envoi_data                     <= '0';  
                    s_plateau                      <= (others =>'0');
                    buffer_plateau                 <= (others =>'0');
                    buff_addr_premier_pixel        <= (others => '0');
                --non utilis� d�sormais mais on garde au cas o�                      
                when etat10 =>
                    -- on indique � la FSM qu'on a fini d'envoyer toutes les donn�es au bloc VGA

                    rst_addr_plateau               <= '0'; 
                    activer_ecriture_vga           <= '0';
                    affectation_cpt_addr_pixel     <= '0';
                    activation_cpt_addr_plateau    <= '0';
                    s_RW_mem                       <= '0';
                    s_activation_memoire           <= '0';  
                    s_fin_affichage                <= '1';
                    envoi_data                     <= '0';
                    s_plateau                      <= (others =>'0');
                    buffer_plateau                 <= (others =>'0');
                    buff_addr_premier_pixel        <= (others => '0');
            end case;    
     end process;
end Behavioral;
